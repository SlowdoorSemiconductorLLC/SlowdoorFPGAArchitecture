module a(b, c, d, e);inout wire [1:0] b;inout wire [1:0] c;inout wire [1:0] d;inout wire [1:0] e;reg [2:0] f;reg [3:0] g;assign b[1] = ( c[0] | d[0] | e[0] ) & ( ( ( ( ( ~ c[1] ) & ( ~ d[1] ) & g[0] ) | ( ( ~ c[1] ) & d[1] & g[1] ) | ( c[1] & ( ~ d[1] ) & g[2] ) | ( c[1] & d[1] & g[3] ) ) & ( ( ~ f[2] ) & f[1] & f[0] ) ) | ( ( ( ( ~ c[1] ) & ( ~ e[1] ) & g[0] ) | ( ( ~ c[1] ) & e[1] & g[1] ) | ( c[1] & ( ~ e[1] ) & g[2] ) | ( c[1] & e[1] & g[3] ) ) & ( f[2] & ( ~ f[1] ) & ( ~ f[0] ) ) ) | ( ( ( ( ~ d[1] ) & ( ~ e[1] ) & g[0] ) | ( ( ~ d[1] ) & e[1] & g[1] ) | ( d[1] & ( ~ e[1] ) & g[2] ) | ( d[1] & e[1] & g[3] ) ) & ( f[2] & ( ~ f[1] ) & f[0] ) ) );assign b[0] = c[0] | d[0] | ( e[0] );assign c[1] = ( b[0] | d[0] | e[0] ) & ( ( ( ( ( ~ b[1] ) & ( ~ d[1] ) & g[0] ) | ( ( ~ b[1] ) & d[1] & g[1] ) | ( b[1] & ( ~ d[1] ) & g[2] ) | ( b[1] & d[1] & g[3] ) ) & ( ( ~ f[2] ) & ( ~ f[1] ) & f[0] ) ) | ( ( ( ( ~ b[1] ) & ( ~ e[1] ) & g[0] ) | ( ( ~ b[1] ) & e[1] & g[1] ) | ( b[1] & ( ~ e[1] ) & g[2] ) | ( b[1] & e[1] & g[3] ) ) & ( ( ~ f[2] ) & f[1] & ( ~ f[0] ) ) ) | ( ( ( ( ~ d[1] ) & ( ~ e[1] ) & g[0] ) | ( ( ~ d[1] ) & e[1] & g[1] ) | ( d[1] & ( ~ e[1] ) & g[2] ) | ( d[1] & e[1] & g[3] ) ) & ( f[2] & ( ~ f[1] ) & f[0] ) ) );assign c[0] = b[0] | d[0] | ( e[0] );assign d[1] = ( b[0] | c[0] | e[0] ) & ( ( ( ( ( ~ b[1] ) & ( ~ c[1] ) & g[0] ) | ( ( ~ b[1] ) & c[1] & g[1] ) | ( b[1] & ( ~ c[1] ) & g[2] ) | ( b[1] & c[1] & g[3] ) ) & ( ( ~ f[2] ) & ( ~ f[1] ) & ( ~ f[0] ) ) ) | ( ( ( ( ~ b[1] ) & ( ~ e[1] ) & g[0] ) | ( ( ~ b[1] ) & e[1] & g[1] ) | ( b[1] & ( ~ e[1] ) & g[2] ) | ( b[1] & e[1] & g[3] ) ) & ( ( ~ f[2] ) & f[1] & ( ~ f[0] ) ) ) | ( ( ( ( ~ c[1] ) & ( ~ e[1] ) & g[0] ) | ( ( ~ c[1] ) & e[1] & g[1] ) | ( c[1] & ( ~ e[1] ) & g[2] ) | ( c[1] & e[1] & g[3] ) ) & ( f[2] & ( ~ f[1] ) & ( ~ f[0] ) ) ) );assign d[0] = b[0] | c[0] | ( e[0] );assign e[1] = ( b[0] | c[0] | d[0] ) & ( ( ( ( ( ~ b[1] ) & ( ~ c[1] ) & g[0] ) | ( ( ~ b[1] ) & c[1] & g[1] ) | ( b[1] & ( ~ c[1] ) & g[2] ) | ( b[1] & c[1] & g[3] ) ) & ( ( ~ f[2] ) & ( ~ f[1] ) & ( ~ f[0] ) ) ) | ( ( ( ( ~ b[1] ) & ( ~ d[1] ) & g[0] ) | ( ( ~ b[1] ) & d[1] & g[1] ) | ( b[1] & ( ~ d[1] ) & g[2] ) | ( b[1] & d[1] & g[3] ) ) & ( ( ~ f[2] ) & ( ~ f[1] ) & f[0] ) ) | ( ( ( ( ~ c[1] ) & ( ~ d[1] ) & g[0] ) | ( ( ~ c[1] ) & d[1] & g[1] ) | ( c[1] & ( ~ d[1] ) & g[2] ) | ( c[1] & d[1] & g[3] ) ) & ( ( ~ f[2] ) & f[1] & f[0] ) ) );assign e[0] = b[0] | c[0] | ( d[0] );endmodule
